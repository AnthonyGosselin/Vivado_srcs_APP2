---------------------------------------------------------------------------------------------
--    sig_fct_1.vhd   (temporaire)
---------------------------------------------------------------------------------------------
---------------------------------------------------------------------------------------------
--    Universit� de Sherbrooke - D�partement de GEGI
--
--    Version         : 5.0
--    Nomenclature    : inspiree de la nomenclature 0.2 GRAMS
--    Date            : 29 janvier 2019
--    Auteur(s)       : 
--    Technologie     : ZYNQ 7000 Zybo Z7-10 (xc7z010clg400-1) 
--    Outils          : vivado 2018.2 64 bits
--
---------------------------------------------------------------------------------------------
--  Description 
--  fonction temporaire, aucun calcul
---------------------------------------------------------------------------------------------
--
---------------------------------------------------------------------------------------------
--   � FAIRE:
--   Voir le guide de la probl�matique
---------------------------------------------------------------------------------------------
--
---------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL; 
USE ieee.numeric_std.ALL;
Library UNISIM;
use UNISIM.vcomponents.all;

---------------------------------------------------------------------------------------------
--      FONCTION DISTORTION DURE
---------------------------------------------------------------------------------------------
entity sig_fct_1 is
    Port (  
    i_ech       : in   std_logic_vector (23 downto 0);
    o_ech_fct   : out  std_logic_vector (23 downto 0)                                    
    );
end sig_fct_1;

---------------------------------------------------------------------------------------------

architecture Behavioral of sig_fct_1 is

---------------------------------------------------------------------------------
-- Signaux
----------------------------------------------------------------------------------
    
    CONSTANT Vs : std_logic_vector(21 downto 0) := "1111111111111111111111";
    
---------------------------------------------------------------------------------------------
--    Description comportementale
---------------------------------------------------------------------------------------------
begin 

    process(i_ech)
    begin
        IF abs(to_integer(signed(i_ech))) < Vs then
            o_ech_fct <= i_ech;
        else
            o_ech_fct <= i_ech(23) & '0' & Vs;
        end if;
    end process;
    
end Behavioral;
